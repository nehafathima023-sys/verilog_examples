`timescale 1ns/1ps

module tb_xnor_gate;

    reg a, b;
    wire y;

    // Instantiate DUT
    xnor_gate dut (
        .a(a),
        .b(b),
        .y(y)
    );

    initial begin
        $monitor("Time=%0t | a=%b b=%b -> y=%b", $time, a, b, y);

        a = 0; b = 0; #10;
        a = 0; b = 1; #10;
        a = 1; b = 0; #10;
        a = 1; b = 1; #10;

        $finish;
    end

endmodule
module xnor_gate (
    input  wire a,
    input  wire b,
    output wire y
);

assign y = ~(a ^ b);

endmodule